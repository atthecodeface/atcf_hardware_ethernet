/** @copyright (C) 2019,  Gavin J Stark.  All rights reserved.
 *
 * @copyright
 *    Licensed under the Apache License, Version 2.0 (the "License");
 *    you may not use this file except in compliance with the License.
 *    You may obtain a copy of the License at
 *     http://www.apache.org/licenses/LICENSE-2.0.
 *   Unless required by applicable law or agreed to in writing, software
 *   distributed under the License is distributed on an "AS IS" BASIS,
 *   WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 *   See the License for the specific language governing permissions and
 *   limitations under the License.
 *
 * @file   tb_8b10b.cdl
 * @brief  Testbench for 8b10b encoder and decoder
 *
 */
/*a Includes */
include "encoding.h"
include "encoders.h"

/*a Module */
module tb_8b10b( clock clk,
                 input bit reset_n,
                 input t_8b10b_symbol     dec_symbol,
                 input t_8b10b_enc_data   enc_data,
                 output t_8b10b_dec_data  dec_data,
                 output t_8b10b_symbol    enc_symbol
)
{
    /*b Nets */
    default clock clk;
    default reset active_low reset_n;
    net t_8b10b_dec_data  dec_data_int ;
    net t_8b10b_symbol    enc_symbol_int;
    clocked t_8b10b_dec_data  dec_data   = {*=0} ;
    clocked t_8b10b_symbol    enc_symbol = {*=0} ;

    /*b Instantiations */
    instantiations: {
        encode_8b10b enc( enc_data <= enc_data,
                          symbol => enc_symbol_int );
        decode_8b10b dec( symbol <= dec_symbol,
                          dec_data => dec_data_int);
        enc_symbol <= enc_symbol_int;
        dec_data <= dec_data_int;

        /*b All done */
    }

    /*b All done */
}

